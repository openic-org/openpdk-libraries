** sch_path: /home/designer/shared/amaru/analog/sg13g2_io/sg13g2_Clamp_N20N0D.sch
.subckt sg13g2_Clamp_N20N0D iovss pad[9] pad[8] pad[7] pad[6] pad[5] pad[4] pad[3] pad[2] pad[1] pad[0] sub
*.PININFO iovss:B pad[9:0]:B sub:B
R1 iovss sub ptap1 A=55.7736p P=328.08u
M1 pad[0] net1 iovss sub sg13_hv_nmos w=8.8u l=0.6u ng=2 m=1
M2 pad[1] net1 iovss sub sg13_hv_nmos w=8.8u l=0.6u ng=2 m=1
M3 pad[2] net1 iovss sub sg13_hv_nmos w=8.8u l=0.6u ng=2 m=1
M4 pad[3] net1 iovss sub sg13_hv_nmos w=8.8u l=0.6u ng=2 m=1
M5 pad[4] net1 iovss sub sg13_hv_nmos w=8.8u l=0.6u ng=2 m=1
M6 pad[5] net1 iovss sub sg13_hv_nmos w=8.8u l=0.6u ng=2 m=1
M7 pad[6] net1 iovss sub sg13_hv_nmos w=8.8u l=0.6u ng=2 m=1
M8 pad[7] net1 iovss sub sg13_hv_nmos w=8.8u l=0.6u ng=2 m=1
M9 pad[8] net1 iovss sub sg13_hv_nmos w=8.8u l=0.6u ng=2 m=1
M10 pad[9] net1 iovss sub sg13_hv_nmos w=8.8u l=0.6u ng=2 m=1
R2 net1 iovss rppd w=0.5e-6 l=3.54e-6 m=1 b=0
.ends
