** sch_path: /home/designer/shared/amaru/analog/sg13g2_io/sg13g2_GateLevelUpInv.sch
.subckt sg13g2_GateLevelUpInv iovdd vss core pgate vdd sub ngate
*.PININFO iovdd:B vss:B pgate:B core:B vdd:B sub:B ngate:B
x1 iovdd vss core pgate vdd sub sg13g2_LevelUpInv_noptap
x2 iovdd vss core ngate vdd sub sg13g2_LevelUpInv_noptap
R1 vss sub ptap1 A=2.106p P=14.64u
.ends

* expanding   symbol:  sg13g2_LevelUpInv_noptap.sym # of pins=6
** sym_path: /home/designer/shared/amaru/analog/sg13g2_io/sg13g2_LevelUpInv_noptap.sym
** sch_path: /home/designer/shared/amaru/analog/sg13g2_io/sg13g2_LevelUpInv_noptap.sch
.subckt sg13g2_LevelUpInv_noptap iovdd vss in out vdd sub
*.PININFO iovdd:B vss:B out:B in:B vdd:B sub:B
M1 net1 in vss sub sg13_hv_nmos w=1.9u l=0.45u ng=1 m=1
M3 net1 net2 iovdd iovdd sg13_hv_pmos w=0.3u l=0.45u ng=1 m=1
M4 net2 net1 iovdd iovdd sg13_hv_pmos w=0.3u l=0.45u ng=1 m=1
M5 out net2 iovdd iovdd sg13_hv_pmos w=3.9u l=0.45u ng=1 m=1
M2 net2 net3 vss sub sg13_hv_nmos w=1.9u l=0.45u ng=1 m=1
M6 out net2 vss sub sg13_hv_nmos w=1.9u l=0.45u ng=1 m=1
M7 net3 in vss sub sg13_lv_nmos w=2.75u l=0.13u ng=1 m=1
M8 net3 in vdd vdd sg13_lv_pmos w=4.75u l=0.13u ng=1 m=1
.ends

