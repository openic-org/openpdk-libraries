* Extracted by KLayout with SG13G2 LVS runset on : 20/02/2026 17:22

.SUBCKT sg13g2_Filler1000 iovss iovss$1 iovss$2 vss
R$1 \$1 vss ptap1 A=1.368p P=9.72u
R$2 \$1 iovss$2 ptap1 A=110.475p P=58.1u
R$3 \$1 iovss$1 ptap1 A=108.27p P=57.12u
R$4 \$1 iovss ptap1 A=110.52p P=58.12u
.ENDS sg13g2_Filler1000
