* Extracted by KLayout with SG13G2 LVS runset on : 20/02/2026 17:24

.SUBCKT sg13g2_Filler2000 iovss iovss$1 iovss$2 vss
R$1 \$1 vss ptap1 A=2.85p P=19.6u
R$2 \$1 iovss$2 ptap1 A=233.225p P=68.1u
R$3 \$1 iovss$1 ptap1 A=228.57p P=67.12u
R$4 \$1 iovss ptap1 A=233.32p P=68.12u
.ENDS sg13g2_Filler2000
