** sch_path: /home/designer/shared/amaru/analog/sg13g2_io/sg13g2_IOPadIn.sch
.subckt sg13g2_IOPadIn vss vdd sub iovss iovdd iovss1 pad p2c
*.PININFO iovdd:B vss:B vdd:B sub:B iovss:B iovss1:B pad:B p2c:B
R2 vss sub ptap1 A=24p P=160.6u
R1 iovss1 sub ptap1 A=5416.1304p P=746.28u
x4 iovdd iovss1 pad p2c vdd vss sub sg13g2_LevelDown_noptap
x2 iovdd sub pad pad sub sg13g2_DCPDiode_noptap
x1 pad iovss pad iovdd sub sg13g2_DCNDiode
.ends

* expanding   symbol:  sg13g2_LevelDown_noptap.sym # of pins=7
** sym_path: /home/designer/shared/amaru/analog/sg13g2_io/sg13g2_LevelDown_noptap.sym
** sch_path: /home/designer/shared/amaru/analog/sg13g2_io/sg13g2_LevelDown_noptap.sch
.subckt sg13g2_LevelDown_noptap iovdd iovss pad core vdd vss sub
*.PININFO iovdd:B vss:B core:B pad:B vdd:B iovss:B sub:B
M5 net2 net1 vdd vdd sg13_hv_pmos w=4.65u l=0.45u ng=1 m=1
M6 net2 net1 vss sub sg13_hv_nmos w=2.65u l=0.45u ng=1 m=1
M7 core net2 vss sub sg13_lv_nmos w=2.75u l=0.13u ng=1 m=1
M8 core net2 vdd vdd sg13_lv_pmos w=4.75u l=0.13u ng=1 m=1
x1 net1 iovdd iovss pad sub sg13g2_SecondaryProtection_noptap
.ends


* expanding   symbol:  sg13g2_DCPDiode_noptap.sym # of pins=5
** sym_path: /home/designer/shared/amaru/analog/sg13g2_io/sg13g2_DCPDiode_noptap.sym
** sch_path: /home/designer/shared/amaru/analog/sg13g2_io/sg13g2_DCPDiode_noptap.sch
.subckt sg13g2_DCPDiode_noptap cathode guard anode1 anode2 sub
*.PININFO anode2:B cathode:B guard:B anode1:B sub:B
D1 anode1 cathode dpantenna l=27.78u w=1.26u
D2 anode2 cathode dpantenna l=27.78u w=1.26u
.ends


* expanding   symbol:  sg13g2_DCNDiode.sym # of pins=5
** sym_path: /home/designer/shared/amaru/analog/sg13g2_io/sg13g2_DCNDiode.sym
** sch_path: /home/designer/shared/amaru/analog/sg13g2_io/sg13g2_DCNDiode.sch
.subckt sg13g2_DCNDiode cathode1 anode cathode2 guard sub
*.PININFO cathode2:B guard:B anode:B cathode1:B sub:B
R1 anode sub ptap1 A=141.2964p P=221.76u
D1 sub cathode1 dantenna l=27.78u w=1.26u
* noconn guard
D2 sub cathode2 dantenna l=27.78u w=1.26u
.ends


* expanding   symbol:  sg13g2_SecondaryProtection_noptap.sym # of pins=5
** sym_path: /home/designer/shared/amaru/analog/sg13g2_io/sg13g2_SecondaryProtection_noptap.sym
** sch_path: /home/designer/shared/amaru/analog/sg13g2_io/sg13g2_SecondaryProtection_noptap.sch
.subckt sg13g2_SecondaryProtection_noptap core iovdd iovss pad sub
*.PININFO iovss:B core:B pad:B iovdd:B sub:B
D1 core iovdd dpantenna l=4.98u w=0.64u
R2 core pad rppd w=1e-6 l=2e-6 m=1 b=0
D2 sub core dantenna l=3.1u w=0.64u
.ends

