** sch_path: /home/designer/shared/amaru/analog/sg13g2_io/sg13g2_Clamp_N8N8D.sch
.subckt sg13g2_Clamp_N8N8D gate iovss pad[3] pad[2] pad[1] pad[0] sub
*.PININFO iovss:B gate:B pad[3:0]:B sub:B
R1 iovss sub ptap1 A=55.7736p P=328.08u
D1 sub gate dantenna l=0.78u w=0.78u
M1 pad[0] gate iovss sub sg13_hv_nmos w=8.8u l=0.6u ng=2 m=1
M2 pad[1] gate iovss sub sg13_hv_nmos w=8.8u l=0.6u ng=2 m=1
M3 pad[2] gate iovss sub sg13_hv_nmos w=8.8u l=0.6u ng=2 m=1
M4 pad[3] gate iovss sub sg13_hv_nmos w=8.8u l=0.6u ng=2 m=1
.ends
