* Extracted by KLayout with SG13G2 LVS runset on : 20/02/2026 17:58

.SUBCKT sg13g2_IOPadAnalog pad iovss iovdd iovdd$1 vss padres
X$1 \$1 iovss padres pad iovdd$1 sg13g2_SecondaryProtection
X$2 iovdd pad pad pad pad pad pad pad pad pad pad sg13g2_Clamp_P20N0D_noptap
X$3 iovdd pad pad sg13g2_DCPDiode_noptap
X$4 \$1 iovss pad pad pad pad pad pad pad pad pad pad sg13g2_Clamp_N20N0D
X$5 \$1 iovss pad pad sg13g2_DCNDiode
R$1 \$1 iovss ptap1 A=4373.9448p P=1112.3u
R$2 \$1 vss ptap1 A=23.85p P=159.6u
.ENDS sg13g2_IOPadAnalog

.SUBCKT sg13g2_SecondaryProtection \$1 iovss core pad iovdd
D$1 \$1 core dantenna A=1.984p P=7.48u m=1
D$2 core iovdd dpantenna A=3.1872p P=11.24u m=1
R$3 pad core rppd w=1u l=2u ps=0 b=0 m=1
R$4 \$1 iovss ptap1 A=9.0304p P=53.12u
.ENDS sg13g2_SecondaryProtection

.SUBCKT sg13g2_DCPDiode_noptap cathode anode anode$1
D$1 anode$1 cathode dpantenna A=35.0028p P=58.08u m=1
D$2 anode cathode dpantenna A=35.0028p P=58.08u m=1
.ENDS sg13g2_DCPDiode_noptap

.SUBCKT sg13g2_DCNDiode \$2 anode cathode cathode$1
D$1 \$2 cathode$1 dantenna A=35.0028p P=58.08u m=1
D$2 \$2 cathode dantenna A=35.0028p P=58.08u m=1
R$3 \$2 anode ptap1 A=141.2964p P=221.76u
.ENDS sg13g2_DCNDiode

.SUBCKT sg13g2_Clamp_P20N0D_noptap iovdd pad pad$1 pad$2 pad$3 pad$4 pad$5
+ pad$6 pad$7 pad$8 pad$9
M$1 iovdd \$5 pad iovdd sg13_hv_pmos L=0.6u W=26.64u AS=14.1192p AD=12.1212p
+ PS=44.2u PD=30.28u
M$3 iovdd \$5 pad$1 iovdd sg13_hv_pmos L=0.6u W=26.64u AS=12.1212p AD=12.1212p
+ PS=30.28u PD=30.28u
M$5 iovdd \$5 pad$2 iovdd sg13_hv_pmos L=0.6u W=26.64u AS=12.1212p AD=12.1212p
+ PS=30.28u PD=30.28u
M$7 iovdd \$5 pad$3 iovdd sg13_hv_pmos L=0.6u W=26.64u AS=12.1212p AD=12.1212p
+ PS=30.28u PD=30.28u
M$9 iovdd \$5 pad$4 iovdd sg13_hv_pmos L=0.6u W=26.64u AS=12.1212p AD=12.1212p
+ PS=30.28u PD=30.28u
M$11 iovdd \$5 pad$5 iovdd sg13_hv_pmos L=0.6u W=26.64u AS=12.1212p AD=12.1212p
+ PS=30.28u PD=30.28u
M$13 iovdd \$5 pad$6 iovdd sg13_hv_pmos L=0.6u W=26.64u AS=12.1212p AD=12.1212p
+ PS=30.28u PD=30.28u
M$15 iovdd \$5 pad$7 iovdd sg13_hv_pmos L=0.6u W=26.64u AS=12.1212p AD=12.1212p
+ PS=30.28u PD=30.28u
M$17 iovdd \$5 pad$8 iovdd sg13_hv_pmos L=0.6u W=26.64u AS=12.1212p AD=12.1212p
+ PS=30.28u PD=30.28u
M$19 iovdd \$5 pad$9 iovdd sg13_hv_pmos L=0.6u W=26.64u AS=12.1212p AD=14.1192p
+ PS=30.28u PD=44.2u
R$41 iovdd \$5 rppd w=0.5u l=12.9u ps=0 b=0 m=1
.ENDS sg13g2_Clamp_P20N0D_noptap

.SUBCKT sg13g2_Clamp_N20N0D \$2 iovss pad pad$1 pad$2 pad$3 pad$4 pad$5 pad$6
+ pad$7 pad$8 pad$9
M$1 iovss \$4 pad \$2 sg13_hv_nmos L=0.6u W=8.8u AS=4.664p AD=4.004p PS=15.32u
+ PD=10.62u
M$3 iovss \$4 pad$1 \$2 sg13_hv_nmos L=0.6u W=8.8u AS=4.004p AD=4.004p
+ PS=10.62u PD=10.62u
M$5 iovss \$4 pad$2 \$2 sg13_hv_nmos L=0.6u W=8.8u AS=4.004p AD=4.004p
+ PS=10.62u PD=10.62u
M$7 iovss \$4 pad$3 \$2 sg13_hv_nmos L=0.6u W=8.8u AS=4.004p AD=4.004p
+ PS=10.62u PD=10.62u
M$9 iovss \$4 pad$4 \$2 sg13_hv_nmos L=0.6u W=8.8u AS=4.004p AD=4.004p
+ PS=10.62u PD=10.62u
M$11 iovss \$4 pad$5 \$2 sg13_hv_nmos L=0.6u W=8.8u AS=4.004p AD=4.004p
+ PS=10.62u PD=10.62u
M$13 iovss \$4 pad$6 \$2 sg13_hv_nmos L=0.6u W=8.8u AS=4.004p AD=4.004p
+ PS=10.62u PD=10.62u
M$15 iovss \$4 pad$7 \$2 sg13_hv_nmos L=0.6u W=8.8u AS=4.004p AD=4.004p
+ PS=10.62u PD=10.62u
M$17 iovss \$4 pad$8 \$2 sg13_hv_nmos L=0.6u W=8.8u AS=4.004p AD=4.004p
+ PS=10.62u PD=10.62u
M$19 iovss \$4 pad$9 \$2 sg13_hv_nmos L=0.6u W=8.8u AS=4.004p AD=4.664p
+ PS=10.62u PD=15.32u
R$21 iovss \$4 rppd w=0.5u l=3.54u ps=0 b=0 m=1
R$22 \$2 iovss ptap1 A=55.7736p P=328.08u
.ENDS sg13g2_Clamp_N20N0D
