* Extracted by KLayout with SG13G2 LVS runset on : 20/02/2026 17:39

.SUBCKT sg13g2_io_inv_x1 i nq vdd vss
M$1 vss i nq \$5 sg13_lv_nmos L=0.13u W=3.93u AS=1.3362p AD=1.3362p PS=8.54u
+ PD=8.54u
M$2 vdd i nq vdd sg13_lv_pmos L=0.13u W=4.41u AS=1.4994p AD=1.4994p PS=9.5u
+ PD=9.5u
R$3 \$5 vss ptap1 A=0.624p P=4.76u
.ENDS sg13g2_io_inv_x1
