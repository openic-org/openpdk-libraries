* Extracted by KLayout with SG13G2 LVS runset on : 20/02/2026 16:49

.SUBCKT sg13g2_Clamp_N20N0D iovss pad pad$1 pad$2 pad$3 pad$4 pad$5 pad$6 pad$7
+ pad$8 pad$9
M$1 iovss \$4 pad \$2 sg13_hv_nmos L=0.6u W=8.8u AS=4.664p AD=4.004p PS=15.32u
+ PD=10.62u
M$3 iovss \$4 pad$1 \$2 sg13_hv_nmos L=0.6u W=8.8u AS=4.004p AD=4.004p
+ PS=10.62u PD=10.62u
M$5 iovss \$4 pad$2 \$2 sg13_hv_nmos L=0.6u W=8.8u AS=4.004p AD=4.004p
+ PS=10.62u PD=10.62u
M$7 iovss \$4 pad$3 \$2 sg13_hv_nmos L=0.6u W=8.8u AS=4.004p AD=4.004p
+ PS=10.62u PD=10.62u
M$9 iovss \$4 pad$4 \$2 sg13_hv_nmos L=0.6u W=8.8u AS=4.004p AD=4.004p
+ PS=10.62u PD=10.62u
M$11 iovss \$4 pad$5 \$2 sg13_hv_nmos L=0.6u W=8.8u AS=4.004p AD=4.004p
+ PS=10.62u PD=10.62u
M$13 iovss \$4 pad$6 \$2 sg13_hv_nmos L=0.6u W=8.8u AS=4.004p AD=4.004p
+ PS=10.62u PD=10.62u
M$15 iovss \$4 pad$7 \$2 sg13_hv_nmos L=0.6u W=8.8u AS=4.004p AD=4.004p
+ PS=10.62u PD=10.62u
M$17 iovss \$4 pad$8 \$2 sg13_hv_nmos L=0.6u W=8.8u AS=4.004p AD=4.004p
+ PS=10.62u PD=10.62u
M$19 iovss \$4 pad$9 \$2 sg13_hv_nmos L=0.6u W=8.8u AS=4.004p AD=4.664p
+ PS=10.62u PD=15.32u
R$21 iovss \$4 rppd w=0.5u l=3.54u ps=0 b=0 m=1
R$22 \$2 iovss ptap1 A=55.7736p P=328.08u
.ENDS sg13g2_Clamp_N20N0D
