** sch_path: /home/designer/shared/amaru/analog/sg13g2_io/sg13g2_io_nor2_x1.sch
.subckt sg13g2_io_nor2_x1 vss i0 nq vdd sub i1
*.PININFO vss:B nq:B i0:B vdd:B sub:B i1:B
R1 vss sub ptap1 A=0.657p P=4.98u
M7 nq i0 vss sub sg13_lv_nmos w=3.93u l=0.13u ng=1 m=1
M8 net1 i0 vdd vdd sg13_lv_pmos w=4.41u l=0.13u ng=1 m=1
M1 nq i1 vss sub sg13_lv_nmos w=3.93u l=0.13u ng=1 m=1
M2 nq i1 net1 vdd sg13_lv_pmos w=4.41u l=0.13u ng=1 m=1
.ends
