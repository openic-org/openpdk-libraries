** sch_path: /home/designer/shared/amaru/analog/sg13g2_io/sg13g2_Clamp_P15N15D.sch
.subckt sg13g2_Clamp_P15N15D gate iovdd iovss pad[7] pad[6] pad[5] pad[4] pad[3] pad[2] pad[1] pad[0] sub
*.PININFO iovss:B gate:B iovdd:B pad[7:0]:B sub:B
R1 iovss sub ptap1 A=67.0344p P=394.32u
M1 pad[0] gate iovdd iovdd sg13_hv_pmos w=26.64u l=0.6u ng=4 m=1
D1 gate iovdd dpantenna l=0.78u w=0.78u
M2 pad[1] gate iovdd iovdd sg13_hv_pmos w=26.64u l=0.6u ng=4 m=1
M3 pad[2] gate iovdd iovdd sg13_hv_pmos w=26.64u l=0.6u ng=4 m=1
M4 pad[3] gate iovdd iovdd sg13_hv_pmos w=26.64u l=0.6u ng=4 m=1
M5 pad[4] gate iovdd iovdd sg13_hv_pmos w=26.64u l=0.6u ng=4 m=1
M6 pad[5] gate iovdd iovdd sg13_hv_pmos w=26.64u l=0.6u ng=4 m=1
M7 pad[6] gate iovdd iovdd sg13_hv_pmos w=26.64u l=0.6u ng=4 m=1
M8 pad[7] gate iovdd iovdd sg13_hv_pmos w=13.32u l=0.6u ng=2 m=1
.ends
