* Extracted by KLayout with SG13G2 LVS runset on : 20/02/2026 16:41

.SUBCKT sg13g2_Clamp_N2N2D iovss gate pad
M$1 iovss gate pad \$2 sg13_hv_nmos L=0.6u W=8.8u AS=4.664p AD=4.664p PS=15.32u
+ PD=15.32u
D$3 \$2 gate dantenna A=0.6084p P=3.12u m=1
R$4 \$2 iovss ptap1 A=55.7736p P=328.08u
.ENDS sg13g2_Clamp_N2N2D
