* Extracted by KLayout with SG13G2 LVS runset on : 20/02/2026 17:25

.SUBCKT sg13g2_Filler4000 iovss iovss$1 iovss$2 vss
R$1 \$1 vss ptap1 A=5.85p P=39.6u
R$2 \$1 iovss$2 ptap1 A=478.725p P=88.1u
R$3 \$1 iovss$1 ptap1 A=469.17p P=87.12u
R$4 \$1 iovss ptap1 A=478.92p P=88.12u
.ENDS sg13g2_Filler4000
