* Extracted by KLayout with SG13G2 LVS runset on : 20/02/2026 17:26

.SUBCKT sg13g2_Filler10000 iovss iovss$1 iovss$2 vss
R$1 \$1 vss ptap1 A=14.85p P=99.6u
R$2 \$1 iovss$2 ptap1 A=1215.225p P=148.1u
R$3 \$1 iovss$1 ptap1 A=1190.97p P=147.12u
R$4 \$1 iovss ptap1 A=1215.72p P=148.12u
.ENDS sg13g2_Filler10000
