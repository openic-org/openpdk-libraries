** sch_path: /home/designer/shared/amaru/analog/sg13g2_io/sg13g2_Filler200.sch
.subckt sg13g2_Filler200 iovdd iovss1 vdd iovss2 iovss3 vss sub
*.PININFO iovss1:B iovss2:B iovss3:B vss:B iovdd:B vdd:B sub:B
R3 iovss3 sub ptap1 A=13.7536p P=50.24u
R4 vss sub ptap1 A=0.678p P=5.12u
R1 iovss1 sub ptap1 A=13.748p P=50.22u
R2 iovss2 sub ptap1 A=13.4736p P=49.24u
* noconn iovdd
* noconn vdd
.ends
