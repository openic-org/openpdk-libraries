** sch_path: /home/designer/shared/amaru/analog/sg13g2_io/sg13g2_Filler2000.sch
.subckt sg13g2_Filler2000 iovdd iovss1 vdd iovss2 iovss3 vss sub
*.PININFO iovss1:B iovss2:B iovss3:B vss:B iovdd:B vdd:B sub:B
R3 iovss3 sub ptap1 A=233.225p P=68.1u
R4 vss sub ptap1 A=2.85p P=19.6u
* noconn iovdd
* noconn vdd
R1 iovss1 sub ptap1 A=233.32p P=68.12u
R2 iovss2 sub ptap1 A=228.57p P=67.12u
.ends
