* Extracted by KLayout with SG13G2 LVS runset on : 20/02/2026 17:46

.SUBCKT sg13g2_LevelUp iovdd o i vss vdd
M$1 \$6 i vss \$5 sg13_lv_nmos L=0.13u W=2.75u AS=0.935p AD=0.935p PS=6.18u
+ PD=6.18u
M$2 vss \$4 o \$5 sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.646p PS=4.48u
+ PD=4.48u
M$3 \$3 \$6 vss \$5 sg13_hv_nmos L=0.45u W=1.9u AS=0.646p AD=0.361p PS=4.48u
+ PD=2.28u
M$4 vss i \$4 \$5 sg13_hv_nmos L=0.45u W=1.9u AS=0.361p AD=0.646p PS=2.28u
+ PD=4.48u
M$5 \$6 i vdd vdd sg13_lv_pmos L=0.13u W=4.75u AS=1.615p AD=1.615p PS=10.18u
+ PD=10.18u
M$6 iovdd \$4 o iovdd sg13_hv_pmos L=0.45u W=3.9u AS=1.326p AD=1.326p PS=8.48u
+ PD=8.48u
M$7 \$3 \$4 iovdd iovdd sg13_hv_pmos L=0.45u W=0.3u AS=0.102p AD=0.057p
+ PS=1.28u PD=0.68u
M$8 iovdd \$3 \$4 iovdd sg13_hv_pmos L=0.45u W=0.3u AS=0.057p AD=0.102p
+ PS=0.68u PD=1.28u
R$9 \$5 vss ptap1 A=0.9135p P=6.69u
.ENDS sg13g2_LevelUp
