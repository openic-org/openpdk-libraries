* Extracted by KLayout with SG13G2 LVS runset on : 20/02/2026 17:20

.SUBCKT sg13g2_Filler200 iovss iovss$1 iovss$2 vss
R$1 \$1 vss ptap1 A=0.678p P=5.12u
R$2 \$1 iovss$2 ptap1 A=13.748p P=50.22u
R$3 \$1 iovss$1 ptap1 A=13.4736p P=49.24u
R$4 \$1 iovss ptap1 A=13.7536p P=50.24u
.ENDS sg13g2_Filler200
