** sch_path: /home/designer/shared/amaru/analog/sg13g2_io/sg13g2_Filler1000.sch
.subckt sg13g2_Filler1000 iovdd iovss1 vdd iovss2 iovss3 vss sub
*.PININFO iovss1:B iovss2:B iovss3:B vss:B iovdd:B vdd:B sub:B
R3 iovss3 sub ptap1 A=110.475p P=58.1u
R4 vss sub ptap1 A=1.368p P=9.72u
* noconn iovdd
* noconn vdd
R1 iovss1 sub ptap1 A=110.52p P=58.12u
R2 iovss2 sub ptap1 A=108.27p P=57.12u
.ends
