** sch_path: /home/designer/shared/amaru/analog/sg13g2_io/sg13g2_Filler4000.sch
.subckt sg13g2_Filler4000 iovdd iovss1 vdd iovss2 iovss3 vss sub
*.PININFO iovss1:B iovss2:B iovss3:B vss:B iovdd:B vdd:B sub:B
R3 iovss3 sub ptap1 A=478.725p P=88.1u
R4 vss sub ptap1 A=5.85p P=39.6u
* noconn iovdd
* noconn vdd
R1 iovss1 sub ptap1 A=478.92p P=88.12u
R2 iovss2 sub ptap1 A=469.17p P=87.12u
.ends
