* Extracted by KLayout with SG13G2 LVS runset on : 20/02/2026 17:17

.SUBCKT sg13g2_DCNDiode anode cathode cathode$1
D$1 \$2 cathode$1 dantenna A=35.0028p P=58.08u m=1
D$2 \$2 cathode dantenna A=35.0028p P=58.08u m=1
R$3 \$2 anode ptap1 A=141.2964p P=221.76u
.ENDS sg13g2_DCNDiode
