* Extracted by KLayout with SG13G2 LVS runset on : 20/02/2026 17:21

.SUBCKT sg13g2_Filler400 iovss iovss$1 iovss$2 vss
R$1 \$1 vss ptap1 A=0.672p P=5.08u
R$2 \$1 iovss$2 ptap1 A=38.298p P=52.22u
R$3 \$1 iovss$1 ptap1 A=37.5336p P=51.24u
R$4 \$1 iovss ptap1 A=38.3136p P=52.24u
.ENDS sg13g2_Filler400
