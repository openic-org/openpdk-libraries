** sch_path: /home/designer/shared/amaru/analog/sg13g2_io/sg13g2_RCClampInverter.sch
.subckt sg13g2_RCClampInverter supply iovss in out sub
*.PININFO supply:B iovss:B out:B in:B sub:B
R1 iovss sub ptap1 A=69.122p P=406.6u
M1 iovss in iovss sub sg13_hv_nmos w=126u l=9.5u ng=14 m=1
M2 out in iovss sub sg13_hv_nmos w=108u l=0.5u ng=12 m=1
M3 out in supply supply sg13_hv_pmos w=350u l=0.5u ng=50 m=1
.ends
