* Extracted by KLayout with SG13G2 LVS runset on : 20/02/2026 17:50

.SUBCKT sg13g2_RCClampInverter iovss in out supply
M$1 iovss in iovss \$1 sg13_hv_nmos L=9.5u W=126u AS=26.64p AD=23.94p
+ PS=149.92u PD=131.32u
M$8 iovss in out \$1 sg13_hv_nmos L=0.5u W=108u AS=20.52p AD=23.22p PS=112.56u
+ PD=131.16u
M$27 supply in out supply sg13_hv_pmos L=0.5u W=350u AS=67.55p AD=67.55p
+ PS=376.3u PD=376.3u
R$77 \$1 iovss ptap1 A=69.122p P=406.6u
.ENDS sg13g2_RCClampInverter
